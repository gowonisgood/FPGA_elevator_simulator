/***********************
*
* Jong-gyu Park
* pjk5401@gmail.com
* 2016/09/02
*
***********************/

module PNU_NOT(i1, o1);
    input i1;
    output o1;
    assign o1=~i1;
endmodule