/***********************
*
* Jong-gyu Park
* pjk5401@gmail.com
* 2016/09/02
*
***********************/

module PNU_AND2(i1, i2, o1);
    input i1, i2;
    output o1;
    assign o1 = i1 & i2;
endmodule